module load_size(

);