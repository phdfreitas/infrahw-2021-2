module store_control(

);